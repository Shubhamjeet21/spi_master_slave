`timescale 1ns / 1ps
package spi_pkg;

  `include "transaction.sv"
  `include "generator.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "environment.sv"

endpackage

